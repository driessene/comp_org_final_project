module ControlUnit ();

endmodule
